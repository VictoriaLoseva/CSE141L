lw $readu
inc
lw $readl
inc
cpy $writeU, $readU
sw $readu 30
inc
cpy $writeL, $readL
sw $readl 30
inc
